`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:56:42 09/25/2014 
// Design Name: 
// Module Name:    q_gen 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module q_gen
	
	
	(
		
	 );

always @ * begin
	if(~nRST) begin
		
	end else begin
	
	end

end

endmodule
